// file: forwarding_unit.v

module forward_unit(
	output wire [1:0] ALU_port1_mux_sel, ALU_port2_mux_sel);
	
	

endmodule